parameter len = 16,  
p = 65521,
g = 373,
q = p - 1